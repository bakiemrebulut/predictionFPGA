
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.types.all;



entity ann is
port 
	(
		clk : in std_logic;
		output : out std_LOGIC;
		reset : in std_LOGIC;
		frame : in img;
		done	: out std_logic
	);

end entity;

architecture rtl of ann is
signal layer : layerarray := ((others=> (others=>'0')));
signal outputSum : std_LOGIC_VECTOR(17 downto 0):=(others=>'0');
signal outputSignal : std_logic:='0';
signal state : std_logic_vector(1 downto 0):="00";	
signal weight :  weightType;
begin 
--oSum<=outputSum(8 downto 0);
output<=outputSignal;
weight <=("000000010101100", "000000100111110", "000000101110001", "000000101011011", "000000101001010", "000000100010000", "000000101111011", "000000101001101", "000000101111001", "000000100010000", "000000011101011", "000000100101110", "000000100110111", "000000010100010", "000000100011011", "000000101100001", "000000010001011", "000000100011110", "000000011110001", "000000100101110", "000000011001101", "000000010101010", "000000010101101", "000000010000111", "000000011100100", "000000011111001", "000000011010100", "000000010010000", "000000101000000", "000000010011111", "000000011010011", "000000101001011", "000000010100111", "000000101011001", "000000011111001", "000000011110001", "000000100100000", "000000011010010", "000000000000000", "000000010011010", "000000011010110", "000000100101011", "000000010011011", "000000010000011", "000000101010001", "000000010101011", "000000100110100", "000000100101010", "000000100101000", "000000100001100", "000000011001100", "000000010100100", "000000010000000", "000000010010010", "000000101100000", "000000101010010", "000000010101101", "000000101000100", "000000100001100", "000000101100110", "000000100110010", "000000100001011", "000000010001000", "000000100001110", "000000011011110", "000000011001000", "000000101010111", "000000101010101", "000000100010010", "000000100101111", "000000011000101", "000000101100010", "000000011101000", "000000101000001", "000000101000110", "000000010010011", "000000011000000", "000000011010111", "000000010001100", "000000101100101", "000000010100101", "000000010110010", "000000011011011", "000000100001101", "000000101101010", "000000100100001", "000000100010000", "000000101000011", "000000100110011", "000000100111111", "000000010111000", "000000100100010", "000000100111010", "000000010101101", "000000000000000", "000000010011110", "000000101110000", "000000010100111", "000000101011011", "000000101100010", "000000011110100", "000000010001011", "000000011111110", "000000011011110", "000000100011100", "000000011010111", "000000010110001", "000000101011001", "000000101101011", "000000011001111", "000000011010100", "000000100010110", "000000100001000", "000000101001110", "000000010011110", "000000101101110", "000000101110110", "000000010001011", "000000011101011", "000000010011100", "000000010010001", "000000011000010", "000000101111110", "000000011011101", "000000100010101", "000000100001000", "000000011111111", "000000010001100", "000000010011100", "000000010000110", "000000100110110", "000000011110100", "000000010011010", "000000100100010", "000000100010101", "000000010110111", "000000100101011", "000000010001110", "000000100100100", "000000010011011", "000000100111111", "000000101010011", "000000101100011", "000000011111011", "000000100100001", "000000101010101", "000000100110111", "000000101010110", "000000101101000", "000000101100011", "000000011010000", "000000011001100", "000000101101100", "000000101100100", "000000010011001", "000000101100110", "000000010010000", "000000101101100", "000000010100110", "000000010001011", "000000100000000", "000000101101110", "000000100010001", "000000101000010", "000000100001010", "000000010110110", "000000010011001", "000000100110111", "000000101111010", "000000011101010", "000000100101011", "000000010111001", "000000011111101", "000000010100001", "000000100111110", "000000101001110", "000000101000101", "000000010000101", "000000100010001", "000000010111010", "000000100000110", "000000010111101", "000000100100110", "000000011110100", "000000010001001", "000000101001010", "000000011001111", "000000011111100", "000000100010000", "000000010001101", "000000101110001", "000000101000111", "000000100001011", "000000010101110", "000000100100110", "000000010011101", "000000100110000", "000000101010001", "000000010111111", "000000100100011", "000000101100110", "000000100010101", "000000010010110", "000000101010110", "000000100000010", "000000011001111", "000000101111000", "000000101011101", "000000010011011", "000000100110000", "000000101110010", "000000010010101", "000000100111010", "000000101001010", "000000101000110", "000000100100111", "000000011101010", "000000100101010", "000000011011101", "000000100001101", "000000010110110", "000000100100101", "000000010100111", "000000100101110", "000000100111010", "000000011111011", "000000101011001", "000000011011010", "000000100000111", "000000100011100", "000000101000101", "000000010011100", "000000101110100", "000000101000010", "000000010011110", "000000011011100", "000000010101101", "000000101000010", "000000010111110", "000000100011111", "000000011111010", "000000101011111", "000000101111110", "000000101010101", "000000100101011", "000000101100100", "000000000000000", "000000010001001", "000000000000000", "000000101000111", "000000000000000", "000000010001100", "000000000000000", "000000101011000", "000000000000000", "000000101110111", "000000010010001", "000000010101011", "000000101100100", "000000010000110", "000000100111101", "000000011111101", "000000100111000", "000000011011011", "000000100010100", "000000010000101", "000000101111010", "000000011100101", "000000101110101", "000000100010000", "000000101010111", "000000101101001", "000000010000110", "000000011111000", "000000100111101", "000000010010100", "000000011100110", "000000100101011", "000000100111110", "000000101110000", "000000100111101", "000000011101000", "000000011001100", "000000010110000", "000000010101000", "000000010100001", "000000101010100", "000000100001011", "000000010010010", "000000101010011", "000000011111000", "000000000000000", "000000101101011", "000000000010000", "000000011100110", "000000000000000", "000000100011010", "000000000000000", "000000101100101", "000000000000000", "000000000101110", "000000100001011", "100001011001001", "000001000000101", "100010010100011", "000001101100100", "100010011001000", "000001100010001", "100010010010101", "000001011000101", "100010000000000", "000001011101101", "100001001101001", "000000110110000", "000000000111101", "000000101000110", "000000010000110", "000000000000000", "000000100011101", "000000000000000", "000000100110010", "000000000000000", "000000011011101", "000000000000101", "000000011001001", "000000010001001", "000000100001100", "000000101000101", "000000100110001", "000000101011000", "000000101000100", "000000101010111", "000000011100100", "000000100111001", "000000100111101", "000000010110010", "000000100110101", "000000010110001", "000000100111101", "000000101011100", "000000011000001", "000000100100111", "000000011110010", "000000011110011", "000000101101011", "000000010100010", "000000100110100", "000000000010001", "000000110000111", "000000001000000", "000001000110001", "000000001111111", "000000111011011", "000000001010110", "100001010011001", "000001000011001", "100001110111000", "000001000101010", "100000111001101", "000000111111000", "100000100101010", "000000011110100", "100000100101011", "000000100010000", "100000101011011", "000000101100110", "100000111001000", "000000111001001", "100001100100110", "000001000101010", "100001111001100", "000001100000101", "100001000111100", "000000111010111", "000001000111011", "000000001010101", "000000110001100", "000000001100111", "000001000010110", "000000001000111", "000000100011010", "000000000001111", "000000010110000", "000000011001001", "000000100101001", "000000101100000", "000000101100001", "000000010011100", "000000011000011", "000000010101110", "000000011100000", "000000011110000", "000000101001110", "000000011101101", "000000101110001", "000000100000011", "000000011011111", "000000100000100", "000000010110110", "000000100000001", "000000101001101", "000000101100011", "000000011000001", "000000000000000", "000001000111110", "000000001101110", "000000001010001", "000000101001001", "100001111100011", "000001010001100", "100000110101110", "000000111110100", "000000011100011", "000000000000000", "000000011101110", "000000000000000", "000001000100001", "000000001011001", "000001000111010", "000000001101001", "000000111011000", "000000001110111", "000001000101001", "000000001011000", "000000011101011", "000000000000000", "000000011001001", "000000101111001", "100001011011110", "000001010111101", "100001110011011", "000001010011110", "000000001000110", "000000000000000", "000000110011011", "000000001011011", "000000101000001", "000000000000000", "000000010011001", "000000000000000", "000000011000001", "000000011111000", "000000011100010", "000000010000010", "000000100110011", "000000100001000", "000000101101001", "000000101010100", "000000100011001", "000000010010001", "000000010001000", "000000010001101", "000000010011000", "000000010111000", "000000011011101", "000000010101110", "000000101011100", "000000010011101", "000000101011110", "000000000000000", "000000110101000", "000000000100110", "100010000011101", "000001011111110", "100000110110100", "000000110011000", "000000011001101", "000000011101010", "000000110010100", "000000000001111", "000001000000101", "000000000100010", "000001000110001", "000000010000100", "000001001010000", "000000010100111", "000001000111101", "000000001111100", "000001011001111", "000000010010101", "000000111101110", "000000001010110", "000000100001100", "000000000010000", "000000001101010", "000000101000011", "100001010110001", "000000111001001", "100001110100010", "000001011011101", "000000110001001", "000000000110000", "000000010110111", "000000000000000", "000000010111101", "000000000000000", "000000100100101", "000000100000101", "000000011010000", "000000010000100", "000000100111111", "000000100010000", "000000101011101", "000000100000011", "000000101010101", "000000101110011", "000000011001000", "000000010001001", "000000011110010", "000000100001010", "000000100011011", "000000010110010", "000000101001100", "000000101111111", "000000010110011", "000000000000000", "100001100000011", "000000111011000", "100000101100001", "000000111010101", "000000011110010", "000000100100011", "000000101100011", "000000000000000", "000000110100011", "000000000010110", "000000011100100", "000000000010110", "000000110000010", "000000001011100", "000001000101111", "000000010011110", "000001001100100", "000000010100001", "000000110110011", "000000001010010", "000000111010011", "000000000111101", "000000101100000", "000000000010011", "000000010110111", "000000000000000", "000000010011100", "000000110010111", "100001011100011", "000001010000001", "100001000011011", "000000110100001", "000000100010111", "000000000000000", "000000101110100", "000000101011100", "000000101110000", "000000011110101", "000000011010110", "000000101110100", "000000010000110", "000000100001101", "000000010011111", "000000100101100", "000000100000111", "000000100001110", "000000100010000", "000000011110000", "000000101111011", "000000011101011", "000000011111001", "000000011111010", "000000100010111", "000000100010010", "000000010010110", "000000011111001", "100001110001111", "000001000111100", "000000010101100", "000000000001010", "000000101010010", "000000000011000", "000000111000110", "000000000000000", "000000011001110", "000000000010110", "000000101110011", "000000000101111", "000001001100111", "000000001100000", "000000111110101", "000000000101011", "000001000100010", "000000000011111", "000001000111010", "000000001011101", "000001000001111", "000000000110011", "000000011111111", "000000000010110", "000000100010100", "000000000000000", "000000100001000", "000000000001001", "000000000000000", "000000000001100", "100001111110010", "000001011010011", "000000001001011", "000000010110110", "000000100100100", "000000010100001", "000000100101011", "000000011011101", "000000011010111", "000000100111000", "000000010011101", "000000011111101", "000000011110100", "000000101111001", "000000010000110", "000000100101111", "000000011001100", "000000011000100", "000000100100100", "000000100000011", "000000100010111", "000000100101000", "000000010100100", "000000010100110", "100001101101110", "000001001111110", "100000100110011", "000000100000101", "000000100001001", "000000000000000", "000000111100011", "000000000011001", "000000011011100", "000000000011010", "000000111001001", "000000000101100", "000001000111010", "000000001101000", "000000100010001", "000000000010100", "000000101110100", "000000000000000", "000000010011000", "000000000000000", "000000111001101", "000000000101110", "000001000100100", "000000000110101", "000000100100001", "000000000111101", "000000100100001", "000000000010110", "000000111100001", "000000000111111", "000000011110001", "000000000010010", "100001010101100", "000001001100110", "100001011011110", "000001000011110", "000000010001000", "000000011000111", "000000010111000", "000000100001011", "000000010110101", "000000010000111", "000000101111001", "000000011110111", "000000010000010", "000000101100111", "000000010011101", "000000101100101", "000000010101111", "000000011001100", "000000101111110", "000000101011101", "000000011001101", "000000011101100", "000000000000000", "000000010101011", "100010011010101", "000001011000000", "100000100100010", "000000110110110", "000000110110000", "000000001011000", "000001001011101", "000000001010011", "000001000101100", "000000001000110", "000000111100111", "000000001011101", "000000101100000", "000000000010100", "000000100110011", "000000000000000", "000000100111100", "000000011110010", "000000100000111", "000000101110111", "000000010111010", "000000000000000", "000000111100000", "000000000011100", "000000111110010", "000000001110101", "000000100100000", "000000000101110", "000000110001100", "000000001101000", "000000110110000", "000000001101000", "100000101111111", "000001000001101", "100010001101100", "000001011010110", "000000000000000", "000000010110001", "000000100110111", "000000010100101", "000000010101011", "000000100001000", "000000101000110", "000000011000101", "000000101101011", "000000100100101", "000000011001101", "000000100000011", "000000100000111", "000000101100001", "000000011111100", "000000101010100", "000000100010110", "000000011000001", "000000000000000", "000000100101101", "100010011101010", "000001110101110", "000000011010100", "000000101101001", "000001001011110", "000000001101000", "000001001110011", "000000001111100", "000001000001001", "000000010100111", "000000100101110", "000000000011001", "000000011100110", "000000000000000", "000000011011111", "000000010111000", "000000011000001", "000000011011011", "000000101100101", "000000101011010", "000000100111111", "000000101110110", "000000100110110", "000000000000000", "000000111100001", "000000001011011", "000001010011110", "000000010001111", "000001000011101", "000000001110000", "000000101111100", "000000001011110", "000000011101110", "000000100010000", "100010011010000", "000001110110010", "000000000000000", "000000101101111", "000000011010101", "000000100001100", "000000011110011", "000000010000101", "000000010010010", "000000010101101", "000000101010110", "000000010000111", "000000011011110", "000000100100100", "000000011011010", "000000101011001", "000000101101111", "000000100011001", "000000010010010", "000000010001000", "000000000000000", "000000100101001", "100010011100100", "000001010111001", "100000100001101", "000000100111101", "000001000011110", "000000001001111", "000000111001000", "000000001111110", "000001010110100", "000000010101001", "000000110011110", "000000000101100", "000000010111110", "000000000000000", "000000101010011", "000000010100101", "000000101001001", "000000100111100", "000000101011011", "000000100101011", "000000101100100", "000000010111100", "000000011111011", "000000000000000", "000000101110011", "000000000101000", "000001101000101", "000000011011111", "000001010000001", "000000001111011", "000000111001000", "000000001010011", "000000011101101", "000000100100111", "100010011110101", "000001110000010", "000000000000000", "000000010001110", "000000101001000", "000000011011110", "000000101010000", "000000101100111", "000000010101011", "000000100110110", "000000011101001", "000000101001010", "000000010011000", "000000101000100", "000000100100010", "000000011100000", "000000100100111", "000000100101110", "000000011000001", "000000100010011", "000000000000000", "000000100010110", "100010001101101", "000001100100111", "100000101011000", "000000111111010", "000000110100001", "000000001011110", "000001000110101", "000000010011111", "000000101111001", "000000000011000", "000000111010000", "000000000010100", "000000011001100", "000000000010011", "000000010001110", "000000000000000", "000000101101010", "000000101010011", "000000101101110", "000000100010101", "000000100101010", "000000000000000", "000000110001011", "000000000010011", "000001000010010", "000000001001000", "000001000110001", "000000001011110", "000001010000110", "000000010100000", "000000111110111", "000000001011110", "100000100110001", "000000100111001", "100010011011011", "000001101011111", "000000000000000", "000000011111100", "000000101100000", "000000010110110", "000000010000011", "000000101011011", "000000010000101", "000000100001100", "000000010010001", "000000010000001", "000000010100000", "000000011010001", "000000100011010", "000000011000111", "000000101110000", "000000101110111", "000000010100101", "000000011000100", "000000101001011", "000000101011110", "100001100100111", "000001010101000", "100000111011101", "000000101011011", "000000111011100", "000000000011101", "000000110101100", "000000001001000", "000000101110101", "000000000100000", "000000101110110", "000000000101000", "000000111110010", "000000000100010", "000000011110111", "000000000010010", "000000011101011", "000000000000000", "000000100010101", "000000000000000", "000000011111000", "000000000010000", "000000110000101", "000000001001001", "000000111011010", "000000000101111", "000000110100100", "000000000010100", "000000111111110", "000000001111100", "000000110001111", "000000000000000", "100000111101111", "000001000111000", "100001101000001", "000001000111111", "000000101000100", "000000101000101", "000000101111101", "000000101111011", "000000101000110", "000000011100000", "000000011001101", "000000011110000", "000000101011011", "000000010100111", "000000101001101", "000000010000000", "000000011111110", "000000101110100", "000000101011100", "000000101000101", "000000011110100", "000000101111100", "000000100000110", "000000100101010", "000000000101010", "000000101101101", "100010000110110", "000001100011010", "000000011100100", "000000000000000", "000000010110111", "000000000000110", "000000100101000", "000000000010010", "000000101010111", "000000000010110", "000000110000010", "000000000100111", "000000110110110", "000000001000011", "000000100001001", "000000000011011", "000000100110111", "000000000100000", "000001000000011", "000000001000111", "000000101010011", "000000000101111", "000000100110101", "000000000010110", "000000011111110", "000000000000000", "000000101010110", "000000000101111", "000000010101010", "000000000010011", "100001101110011", "000001011100011", "000000010010101", "000000100001100", "000000010111101", "000000100101000", "000000101101001", "000000101011010", "000000011001001", "000000100111011", "000000011001001", "000000101000010", "000000100101110", "000000011110110", "000000011001111", "000000101101101", "000000011111101", "000000010000010", "000000010010011", "000000101000010", "000000010000010", "000000011101000", "000000101010000", "000000011101010", "000000011000001", "000000000000000", "100000111100111", "000000111110000", "100001000010010", "000000111001101", "000000001101110", "000000110011001", "000000100100100", "000000000000110", "000000011001110", "000000000000000", "000000011100100", "000000000010110", "000000110100011", "000000000110101", "000000110111011", "000000001111111", "000001000110001", "000000010001101", "000000110000110", "000000000111011", "000000111010000", "000000000011010", "000000100111110", "000000000010010", "000000101110101", "000000000000101", "100000100000100", "000000100001111", "100000101010000", "000000110011100", "100001011010001", "000000111100100", "000000100100001", "000000000000000", "000000100110100", "000000100111101", "000000101110010", "000000010000110", "000000011011001", "000000101101100", "000000011011001", "000000101110101", "000000011100100", "000000101110100", "000000100111101", "000000010001001", "000000100110010", "000000011100100", "000000101010010", "000000101001010", "000000010010010", "000000101000001", "000000100010101", "000000010000000", "000000010101010", "000000000000000", "000001001001010", "000000010011000", "100001110101011", "000001011001000", "100000111110101", "000001001001100", "000000000000000", "000000000101001", "000000100111000", "000000000101011", "000001001001000", "000000001000001", "000000111010110", "000000010000001", "000001001111110", "000000001110110", "000001000001011", "000000010001011", "000001000100110", "000000001111101", "000000101101000", "000000001010001", "000000110110100", "000000000001110", "000000011101000", "000000101011110", "100000110100110", "000000110111001", "100001111001100", "000001001100101", "000000110011001", "000000001010100", "000000010011010", "000000000000000", "000000101000011", "000000101001010", "000000010001001", "000000010100100", "000000101001010", "000000010011010", "000000011010010", "000000101101111", "000000010100001", "000000101001000", "000000101000110", "000000100110000", "000000101101101", "000000101010001", "000000100011110", "000000011111101", "000000011111000", "000000101100110", "000000011101111", "000000100110011", "000000011101011", "000000000000000", "000001000000010", "000000001110100", "000000011011111", "000000000000000", "100001110011010", "000001001100011", "100001001110000", "000000111001010", "000000000011010", "000000000100011", "000000101011001", "000000000101001", "000001010001010", "000000000111101", "000001001010110", "000000001101110", "000001001101011", "000000010000001", "000001001011000", "000000001011101", "000000010011111", "000000000000000", "000000011010000", "000000000000000", "100000110001010", "000000110110010", "100001111001110", "000001001100001", "000000010100011", "000000000000100", "000001011001110", "000000010100000", "000000010100110", "000000000000000", "000000010111011", "000000010011011", "000000010011100", "000000010001000", "000000100010011", "000000011100000", "000000010000101", "000000011011011", "000000101101111", "000000101011101", "000000010001000", "000000010100010", "000000100111110", "000000010111011", "000000010011101", "000000101101001", "000000010101101", "000000101101000", "000000010011101", "000000011010001", "000000110111001", "000000000101000", "000001000111111", "000000000111100", "000000111000111", "000000001111101", "000001001111100", "000000001111011", "100000110111011", "000000110000110", "100001110001110", "000001011000011", "100001010111111", "000001000001101", "100000101111010", "000001000011110", "100000101101001", "000000101100001", "100000100110001", "000000110011000", "100000101111001", "000000100011110", "100001010100010", "000001001011011", "100001111010110", "000001010000001", "100001011000001", "000001001101000", "000000101101111", "000000001000010", "000001000110001", "000000001001100", "000001000110000", "000000001011010", "000000101010110", "000000000000000", "000000010110000", "000000010001010", "000000101010011", "000000010111110", "000000100100111", "000000010011111", "000000010010000", "000000100011010", "000000100010100", "000000100001101", "000000101101011", "000000010000011", "000000101000010", "000000011001011", "000000011000010", "000000010111101", "000000100011001", "000000011010010", "000000010001010", "000000100000100", "000000100000110", "000000000000000", "000000110101111", "000000000011011", "000000101011111", "000000000000000", "000000110000011", "000000000000000", "000000100001100", "000000000000000", "000000000010100", "000000100000100", "100000111100010", "000000111101001", "100001111101001", "000001100111110", "100010000100001", "000001101100101", "100010010101000", "000001101111000", "100010001000001", "000001011001011", "100001010110110", "000001000011100", "000000001101100", "000000010101101", "000000000000000", "000000010110000", "000000011111010", "000000000000000", "000000011111110", "000000000000000", "000000011101010", "000000000010011", "000000100010101", "000000000000000", "000000100001000", "000000101101110", "000000101110111", "000000101001000", "000000010001011", "000000011111001", "000000010111000", "000000010000110", "000000101010111", "000000011111001", "000000100001100", "000000010010111", "000000010000101", "000000011011110", "000000100100010", "000000100001100", "000000101000010", "000000100000110", "000000011011000", "000000010010010", "000000011010010", "000000100100011", "000000011100001", "000000010000100", "000000101101001", "000000011100110", "000000010101100", "000000011101100", "000000100101010", "000000101011101", "000000010010111", "000000101101110", "000000000000000", "000000010011100", "000000000000000", "000000010000111", "000000000000000", "000000101111101", "000000000000000", "000000101110001", "000000000000000", "000000010110101", "000000000000000", "000000010100001", "000000011011111", "000000100110010", "000000101000000", "000000101110110", "000000100011011", "000000011100011", "000000011110110", "000000011001001", "000000100001000", "000000011001110", "000000010101101", "000000101000011", "000000100010000", "000000100001111", "000000011110111", "000000011000111", "000000011100100", "000000101010001", "000000100011110", "000000011110010", "000000010001010", "000000010100001", "000000100111111", "000000101000010", "000000100010010", "000000100100011", "000000010111110", "000000011110111", "000000010111001", "000000011001010", "000000010010000", "000000010110001", "000000011100000", "000000011010010", "000000101111110", "000000100101001", "000000100000010", "000000011111110", "000000100110000", "000000010011101", "000000010101010", "000000011001110", "000000011011100", "000000100110011", "000000011001011", "000000101011111", "000000101101001", "000000100010110", "000000010100010", "000000011001101", "000000101110010", "000000100001010", "000000101000110", "000000011101011", "000000011100101", "000000101011000", "000000010100000", "000000100011110", "000000011111110", "000000100110011", "000000011101101", "000000101111010", "000000010110100", "000000101111110", "000000100111011", "000000101000000", "000000011011110", "000000011000000", "000000011010111", "000000100001100", "000000101110011", "000000100101010", "000000101001101", "000000011110001", "000000010110101", "000000100011000", "000000101000100", "000000011101000", "000000101100000", "000000011110111", "000000010110010", "000000101101100", "000000101111011", "000000101111011", "000000100011110", "000000100001110", "000000100001000", "000000101001010", "000000100110111", "000000010010100", "000000100001000", "000000100001110", "000000101010001", "000000010101110", "000000011000100", "000000010001001", "000000011101100", "000000101000101", "000000011000010", "000000010110101", "000000100010000", "000000010111100", "000000100010000", "000000101100100", "000000101100100", "000000011010110", "000000010101101", "000000011001010", "000000100010011", "000000010000111", "000000101110001", "000000100010110", "000000101011100", "000000011000010", "000000010100101", "000000100110100", "000000010111010", "000000010110010", "000000100001111", "000000010111000", "000000100100000", "000000011010110", "000000010001010", "000000100101011", "000000011010101", "000000010010101", "000000101000010", "000000010110110", "000000010000010", "000000101000100", "000000100110011", "000000101101100", "000000100001101", "000000011110010", "000000101010001", "000000100100111", "000000011011011", "000000011100011", "000000010111101", "000000010010100", "000000101111010", "000000101101001", "000000010100001", "000000010101001", "000000101001000", "000000100001111", "000000010000010", "000000101001011", "000000011101100", "000000010011001", "000000100110111", "000000101001110", "000000010011100", "000000011110100", "000000100011100", "000000010111011", "000000010110000", "000000100011010", "000000101011100", "000000011101111", "000000100111111", "000000010010011", "000000100110101", "000000100101100", "000000100000000", "000000100101100", "000000101110111", "000000101110000", "000000011000000", "000000101100011", "000000010101100", "000000101011010", "000000011001110", "000000011110001", "000000010111011", "000000010111110", "000000101011000", "000000100111100", "000000011111100", "000000101000100", "000000010010000", "000000100001000", "000000101110011", "000000011100110", "000000011111111", "000000010110001", "000000100111100", "000000011001011", "000000101110100", "000000011000011", "000000100010110", "000000011011010", "000000010010111", "000000011010011", "000000010110001", "000000011010000", "000000010110000", "000000100000001", "000000010100101", "000000011100100", "000000101100011", "000000101011001", "000000011010110", "000000011101001", "000000101111111", "000000010010000", "000000010111010", "000000101011100", "000000101110010", "000000100011111", "000000010101110", "000000101111011", "000000010111001", "000000010111110", "000000100110010", "000000101010010", "000000101011101", "000000100110101", "000000010110011", "000000010101000", "000000100001001", "000000010111000", "000000100001100", "000000101110100", "000000101011101", "000000101011100", "000000100101101", "000000100000011", "000000101100111", "000000100101011", "000000101111111", "000000011110101", "000000010000100", "000000100000000", "000000011100000", "000000011010100", "000000100011111", "000000100100100", "000000010001100", "000000010000000", "000000010011111", "000000010100010", "000000011010010", "000000011010100", "000000100011011", "000000010011010", "100011111111001", "000010000000000"); 
process(reset,clk)
variable i : integer range 0 to 784:=0;
	begin 
	if(reset = '1') then
		i:=0;
		state<="00";
		done<='0';
	elsif(rising_edge(clk)) then
		case state is 
			when "00"=>
				if i<=783 then
					layer(0)<=sum1815(x=>layer(0),y=>mulIw1(I=>frame(i),w1=>weight(i*2)));
					layer(1)<=sum1815(x=>layer(1),y=>mulIw1(I=>frame(i),w1=>weight(i*2+1)));
					i:=i+1;
				else	
					layer(0)<=sigmoid18(layer(0));
					layer(1)<=sigmoid18(layer(1));
					state <="01";
				end if;
			when "01"=>
				outputSum<=sum1515(x=>mullw2(	l1=>layer(0),w2=>weight(1568)	),y=>mullw2(l1=>layer(1),w2=>weight(1569)));
				state <="10";
			when "10"=>
			outputSum<=sigmoid18(outputSum);
			state<="11";
			when others=>
			done<='1';
		end case;
	end if;
end process;
outputSignal<=(outputSum(8) or outputSum(7));

end rtl;
