
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.types.all;



entity ann is
port 
	(
		clk : in std_logic;
		output : out std_LOGIC;
		reset : in std_LOGIC;
		oSum : out std_LOGIC_VECTOR(17 downto 0);
		stout : out std_LOGIC_vector(1 downto 0);
		selecttest : in std_logic_vecTOR(1 downto 0):="00";
		testO : out img;
		layerO: out layerarray
		
	);

end entity;

architecture rtl of ann is

signal layer : layerarray := ((others=> (others=>'0')));

signal outputSum : std_LOGIC_VECTOR(17 downto 0):=(others=>'0');


signal outputSignal : std_logic:='0';
signal state : std_logic_vector(1 downto 0):="00";	

signal weight :  weightType;
signal test   :  img;

begin 
stout<=state;
oSum<=outputSum;
output<=outputSignal;
weight <=("000011100110011", "000100100110100", "000010001110000", "000000111010011", "000001111010100", "000010100010010", "000100100101100", "000011011011110", "000011001000111", "000100100110001", "000000000101011", "000011101100001", "000100111100001", "000011011111101", "000000111101011", "000001100010000", "000010011101010", "000001111100010", "000100111101010", "000001111010101", "000011111101001", "000001111011010", "000000010000100", "000000000000000", "100000101010001", "000010101011111", "000000000000000", "000000001000001", "000000000000000", "000000000000000", "000010001111010", "000000000011000", "000000000000000", "000001001010110", "000000001100101", "000010010001101", "000100110111101", "000100111111000", "000000000000000", "000000000000000", "100001110101111", "000000100001000", "100001110101111", "000001001110111", "000000000000000", "000010010001010", "000100000100010", "000000101101000", "000100001111011", "000000101100011", "000000001110111", "000011101000001", "000011001111011", "000010101011011", "000001111010011", "000000100110011", "000100011101110", "000010010001010", "000100100001010", "000010010010011", "000000001101011", "000000000000000", "000000101110101", "000000000000000", "000001111011010", "000000000000000", "000000000000000", "000000000000000", "000000000110010", "000000001010000", "100001010100111", "000000010100001", "100001000101111", "000000110011111", "100010011001110", "000000100101110", "100111011011001", "000001110001101", "100110100101111", "000011010101011", "100011010111110", "000000101000101", "100011110111011", "000001001011000", "100001100100010", "000000011000001", "000110110101110", "000000000000000", "000001111101010", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000000001101000", "100010001100000", "000000100111000", "100001000110110", "000000001000011", "100001001001001", "000000001000011", "000100011111101", "000000000000000", "000010011010110", "000000000000000", "000011101001101", "000000000000000", "000000001011100", "000010111101001", "000000100010111", "000010011101011", "000010011111010", "000001111011010", "000000010110010", "000001100101110", "000100101101100", "000010011101010", "000000101011001", "000000000000000", "100001110001011", "000000011100011", "000000000000000", "000001011011011", "000001000100000", "000000111110011", "000000000000000", "000001001011110", "000000000110101", "000000010001101", "000001110110001", "000000000000000", "000001110001000", "000000000000000", "000001110110101", "000000000000000", "000000000000000", "000001001000110", "000000110001111", "000000000000000", "000000100101011", "000000000000000", "100100001100001", "000000101000111", "101001010100110", "000010010100110", "000010001000111", "000000000000000", "000000101111001", "000000000000000", "000000000000000", "000001000100101", "000000000000000", "000010011101010", "000011000010111", "000000000000000", "000001010000101", "000000000000000", "000000000000000", "000001100111110", "000000101100100", "000000000000000", "000000000110110", "000000000000000", "000011001001100", "000000000011011", "000001010101000", "000011100100100", "000010110000111", "000001100000001", "100001111101110", "000000101001110", "100001001011101", "000010110011101", "000000000000000", "000000000000000", "100010100001101", "000000000000000", "000100010010010", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000000100011001", "000000000000000", "000000000000101", "000000000000000", "100100011111000", "000001000001110", "100100010101001", "000000000000000", "100001001110101", "000000000000000", "100001010100101", "000000000000000", "110000110111111", "000010100011110", "100111100010001", "000000111001100", "100100110010111", "000000110011001", "000000000000000", "100000100010010", "100111010001001", "000100000011100", "000010100111100", "000000000000000", "000010010000011", "000000000000000", "000000000000000", "000000111011111", "000001011100011", "000000000000000", "000000000000000", "000000000000000", "000001111000101", "000000000000000", "000011100011100", "000001000111001", "000001110010001", "000000000000000", "100001111101110", "000001101100110", "000100010010111", "000000010001000", "000000000000000", "000001100000111", "000101001001101", "000000000000000", "001001000010111", "000000011010010", "000000000000000", "000001011011001", "000000001100011", "000000000000000", "000101101101110", "000001001010111", "000000000000000", "000000110000001", "000000000000000", "000000110000000", "100011001000010", "000011010110000", "100000100111000", "000000100010001", "000111000000011", "100000101000111", "000000011011001", "000001011001110", "100111000110001", "000010110001101", "100111110111011", "000000100100100", "100101001110010", "000001010000111", "100100000110010", "000001111100011", "000011010100011", "100001000011001", "000000001101111", "000000000000000", "000001100111000", "000000000000000", "000011011110001", "000000000000000", "000011000101001", "000000000000000", "000111001001001", "100000100111011", "000000000000000", "000000000000000", "000001001100011", "000010001000111", "000001011100110", "000010010001100", "000100001010110", "000000001011101", "000100000110011", "000001011111111", "000000000000000", "000000111100111", "000010010111001", "000000011011110", "000011100010001", "100000100100000", "000010011010101", "000000000000000", "000000010011010", "000000101100100", "000101000001011", "000000000000000", "000111100000000", "000000000000000", "000010000111001", "000000000000000", "000000000000000", "000000000000000", "000000000011010", "000010010101001", "000010100110111", "000000000000000", "100110111011000", "000001001110100", "101000101111011", "000001011000110", "101010001011001", "000011001111011", "100001001100010", "000010101100000", "100000111001011", "000000000000000", "100011011011110", "000001101000110", "000000011111010", "000000001001001", "101000001000110", "000001011011111", "100101101010100", "000000001110011", "000000000010001", "000000000000000", "000011010110101", "000000000000000", "000000011010110", "000000000000000", "000000000000000", "000000000000000", "000100010011100", "000000000000000", "000100100010000", "000001110011110", "000011110101001", "000000000000000", "000100101011100", "000000101000001", "000000000000000", "000001111011110", "000000000000000", "000000111011010", "000100011110010", "100000100011110", "000000000000000", "000000000000000", "000000000001111", "000001101101111", "000000000000000", "000000000000000", "000101001011110", "000000000000000", "101000000011110", "000010100001011", "000011111110100", "000000000000000", "000001011010100", "000000000000000", "100011011011101", "000000010010010", "101100001100010", "000010110001110", "000111110000111", "000000000000000", "100100010111100", "000001000111101", "000000000000000", "000000000000000", "101010100101110", "000100101100111", "000000110100100", "000000000000000", "001000100110111", "100000110010011", "100010011011000", "000001100000110", "010000001001111", "000000000011010", "100111010011110", "000011101111000", "001000001101101", "000000000000000", "000101000001011", "000000000000000", "100001110111001", "000000000111100", "000110111110001", "000000000000000", "000000101100010", "000000000000000", "000000011011010", "000000000000000", "000100000000011", "000010110011010", "000000000000000", "000010000100001", "000000000000000", "000000000000000", "000111001000000", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000000100011111", "000000000100110", "100101111010100", "000000000010000", "000001000001000", "000000000000000", "000011010100110", "000000000000000", "100100101001000", "000001010000011", "000000011001100", "000001110010011", "000011000111110", "000000000000000", "000010011100000", "000001000010110", "100001001000111", "000000000000000", "000000111100010", "000001101111100", "101000101110001", "000100001110011", "100111110000011", "000001100111110", "100000101111101", "000001001000000", "101000111001111", "000011000010101", "101101111110100", "000011010011011", "000000101010100", "000000000000000", "000000000000000", "000000000000000", "000101110111000", "000000000000000", "000000000000000", "000000100111010", "000010011000011", "000000000000000", "000100101010100", "000000000000000", "000100000001110", "000001000001000", "000000010100101", "000100110100010", "000000000000000", "000000000000000", "000000000000000", "000000110100111", "000000000000000", "000000000000000", "000000110100010", "000000000000000", "101000110111011", "000011001111101", "000000000000001", "000000000000000", "100110011100000", "000010000101000", "101100111100100", "000100101011010", "101000100000100", "000000111101001", "100011110110011", "000010111100000", "010000101110111", "000000000000000", "001000000001111", "000000000000000", "001000011100010", "000000000000000", "100111010110111", "000001111011011", "100011101100001", "000001101011011", "000110000111110", "000000000000000", "000000000000000", "000000000000000", "000000010101000", "000000000000000", "000000000000000", "000000000000000", "100110001111001", "000001000011011", "001010011101000", "100001011110100", "100001001011100", "000000000000000", "100011011101010", "000001100100011", "000000000000000", "000000011111100", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000011100011000", "000010010011000", "000001100011100", "000010000111111", "000000000000000", "000000000000010", "000000000000000", "000000000000000", "100111100001001", "000001010111111", "000110001101100", "000000000000111", "000000001100011", "000000000000000", "000011110111000", "000000000000000", "000011010001100", "000000000000000", "101000111110111", "000010010000110", "000101001110101", "000000000000000", "000000000011010", "000001110010111", "001001010011110", "000000000000000", "000101010100010", "000000000000000", "100100101111100", "000011001011001", "000101110001010", "000000000000000", "000000110101100", "000000000000000", "000011111010110", "000000101111110", "101011100111001", "000100010110100", "000000000000000", "000000000000000", "000101111001001", "000000000000000", "000001010000011", "000000000000000", "000110101111110", "000000011100001", "000000000110000", "000000000000000", "100101111101000", "000010100011010", "000000101101111", "000000100111100", "100000100010100", "000000100110110", "000001110001010", "000000000000000", "000100101110010", "000001011011101", "100001001110010", "000010011010110", "100000111010011", "000000000000000", "101000111110010", "000001011111100", "000100110000100", "000000000000000", "000110001000111", "000000001011010", "000101010010101", "000001010110101", "000000000001111", "000000000000000", "000000010111011", "000001011011111", "000011001111101", "000000000000000", "100101010101000", "000010110100000", "100010100011010", "000000000000000", "000000000110110", "000000000000000", "100111110110000", "000010100100010", "000000001110011", "000000000000000", "000010100101001", "000000000000000", "000010011101010", "000000000000000", "001111010010000", "000000011011110", "010010100011100", "000000010110000", "100011100011110", "000010100101001", "100100101110111", "000000101100000", "000000010010110", "000000000000000", "100011010011000", "000001001000100", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "100010001101001", "000000100110011", "100010000011001", "000011100110111", "000000000000000", "000000101100001", "000000000000000", "000000010001100", "000000000011100", "000010011111011", "000000000000000", "000000010110001", "101000101010011", "000001101101100", "100011010011000", "000000011100010", "001100000001011", "000000000000000", "100101000100011", "000001110000111", "100101010001111", "000010010101000", "101010010010010", "000011110011110", "100001010011110", "000001100010101", "000001101011010", "000000000000000", "100100001100001", "000011000011111", "000000000000000", "000000000000000", "000000000000000", "000000110111100", "000000000000000", "000001100001000", "001010111001110", "100010001001001", "001001011100010", "000000000000000", "000000000000000", "000011101110000", "000000000000000", "000001011110011", "010010011111000", "100010110100000", "100001011010001", "000010111110111", "000010000100101", "000000000000000", "100000111100100", "000000000000000", "100101100100110", "000000000000000", "100011000000111", "000000000000000", "000001101110000", "000001011000111", "100011001100010", "000000100011010", "000001010101000", "000000000000000", "000000001101000", "000000010100101", "100010100000011", "000100010001111", "100010100010100", "000001010001010", "100010001110111", "000001000001110", "100010111011001", "000010011011011", "100010000001010", "000001100011010", "000011110100001", "000000000000000", "100001011000010", "000000000000000", "000000011011110", "000000100001011", "000101010001111", "000000000000000", "001011001101111", "000000000000000", "000001010010111", "000000111111011", "000010001101111", "000000000000000", "000000000000000", "000000000000000", "000000111010010", "000000000101011", "000000100010001", "000010101000110", "000110001001111", "000000000000000", "000000000000000", "000000000000000", "000011110011111", "000000000000000", "000000000000000", "000000110000110", "101110111011001", "000011111010011", "000000011011110", "000000000000000", "101010110110010", "000011001010010", "000000001100011", "000000000000000", "100010110010100", "000010000110101", "000010111011000", "000010000101111", "101000001110010", "000100000111110", "000000000000000", "000001010001000", "000000000000000", "000000100001111", "000000010110010", "000001110111111", "100101100110101", "000001101001011", "000000000000000", "000001010110110", "000000000000000", "000000000000000", "000000000000000", "000001011000110", "000000000000000", "000011100100000", "000000000000000", "000000000000000", "000001100010110", "000000000000000", "100001011110110", "000010011000110", "000000000000000", "000000000000000", "000101001001010", "000000000000000", "100010000100001", "000001000001100", "100001010101111", "000001111100001", "000000000000000", "000000000000000", "001010000100010", "000000000000000", "000010101111000", "000000101101111", "100001100010100", "000001111011001", "100101001100001", "000010110110111", "000000000101111", "000010100000000", "000110000111101", "000000000000000", "101001010110111", "000001000101100", "000000111100000", "000000000000000", "001010010110010", "100000111110001", "101001001001010", "000001001110001", "000000000000000", "000011110100101", "100101101111011", "000010011000001", "100011000110111", "000000100101111", "000000011100011", "000000000000000", "100000100101110", "000001010101100", "000000011000000", "000000111011000", "100110100001111", "000011100000100", "100100100000100", "000011001001110", "100011111110101", "000001110110010", "100101010100101", "000010000110101", "000001110110011", "000001001100011", "000101000011100", "000000000000000", "001000101001111", "000000001100000", "001011011011001", "100001100111100", "000000000000000", "000000000000000", "000110101111001", "000000000000000", "110000010010111", "000101100001100", "100111110110000", "000010000101101", "000010100100111", "000000000000000", "000001110000110", "000000000000000", "000111000011101", "000000000000000", "000101000100100", "000001101011011", "001111000101111", "000000000000000", "100111110001011", "000001111011001", "000010010010110", "000000000000000", "100010100101010", "000001010100000", "100010100110111", "000001001001001", "101000011100010", "000001110100001", "000000000000000", "000000000000000", "100011101010101", "000001000011101", "000000000000000", "000000000000000", "000100001111101", "000000000000000", "100001001110010", "000001010001101", "100000111001010", "000000011001011", "101010000001110", "000100010000011", "000000000000000", "000000000000000", "100100101111010", "000101111000111", "000111001110011", "000000000000000", "100110110100100", "000001101010000", "001001101011110", "000000000000000", "000000000000000", "000001001100111", "000110011110100", "000000000000000", "100010010111100", "000000111101010", "000011011011001", "000000000000000", "001011110001100", "000000000000000", "000000000000000", "000000011011011", "000011111001011", "000000000000000", "000100011000110", "000000000000000", "100000100110000", "000011110010010", "001101101111000", "000000000000000", "000100010111011", "000000111001101", "000011010100110", "000000000000000", "100011010100110", "000000001101100", "000000011100001", "000010110010011", "000101111111100", "000000000000000", "000000000000000", "000000000000000", "000010111000110", "000000000000000", "100000101111110", "000000000000000", "000000000000000", "000000000000000", "000010000010101", "000000000000000", "000000000000000", "000000010111111", "100111001110000", "000011110011010", "100110100111101", "000000110101011", "000011100011001", "000000000000000", "100000101111000", "000000000000000", "000110010110011", "000001100110111", "100000100111000", "000010010010000", "000000000000000", "000000001100001", "001010101010010", "000000000000000", "100010101101110", "000001011101100", "000001000100110", "000000000000000", "000000001101101", "000000000000000", "000010100011000", "000000001110110", "001010011010010", "000000000000000", "101011000111101", "000101111100000", "000000000000000", "000010001100100", "001100100001001", "000000000000000", "010011001100001", "000000010001010", "001100010000011", "000000000000000", "000001110001011", "000000000000000", "100010010110011", "000000000000000", "000111111111000", "000000000000000", "100001010001001", "000000001010000", "100001100001111", "000000101000010", "100110100010001", "000100001011101", "100011010100110", "000000001110001", "100010111100111", "000000010010001", "000010001010011", "000000010111111", "100000111001100", "000001101010100", "100111111000100", "000010111000011", "101000000101001", "000100100001101", "000101001010000", "000000000000000", "000001001011001", "000000000000000", "000111100011110", "000000000000000", "100001100011000", "000000111111100", "000000010111100", "000001011011010", "000001000010110", "000000000000000", "100100000100100", "000001100001101", "000010100010100", "000000000000000", "000110111010111", "000000000110000", "000101100111010", "000000000000000", "000000000000000", "000000100011101", "000010010100101", "000000000000000", "000110110111000", "000000000000000", "100001100010011", "000000000000000", "000100000100000", "000000000000000", "001010011001001", "000000000000000", "000000000000000", "000000101100111", "001011100100011", "000000000000000", "000011101111111", "000000000000000", "000000000000001", "000000000000000", "000100001000000", "000000000000000", "101000000011010", "000010011101011", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000001010100100", "000000000000000", "100001001110010", "000000010111111", "100100111111000", "000000110110011", "100001100111100", "000000001001010", "100111101010001", "000011110100001", "000000000000000", "000000111000101", "001101110111100", "100001111011001", "000000000000000", "000010000110011", "100010000101111", "000000001010110", "100010110001010", "000000000000000", "000000000101100", "000000000000000", "100000111000011", "000000000000000", "000000000000000", "000000000000000", "000100110011001", "000000000000000", "100001010100110", "000011110111110", "000011100110001", "000000000000000", "000000000001010", "000001100111011", "100111001101000", "000011001001110", "000100101000011", "000000011000101", "000000000000000", "000000000000000", "100010100010111", "000000011011001", "100001000011010", "000011101101011", "100001101111000", "000000111011110", "000011000001010", "000000000000000", "000000000000000", "000000011011111", "100001110000100", "000000011000000", "000101101010000", "000000000000101", "000000000000000", "000000000000000", "000000010011110", "000000000000000", "000000000000000", "000000000000000", "100000110000110", "000000000000000", "000001001101100", "000000000000000", "000000110000100", "000001010100011", "100110011010110", "000001111000001", "000011110101111", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "101010001100010", "000011110110110", "100001101000110", "000000010011111", "000001011111001", "000000000000000", "100011100100000", "000010001001101", "100000100110111", "000001001000100", "100010101010111", "000001011011110", "101001101010110", "000100001000001", "000000111111011", "000000000000000", "000000110001111", "000000000000000", "000110010011010", "000000000000000", "100011001111110", "000000111000110", "100000100111000", "000000110011001", "101001000111010", "000010111001011", "000000010010001", "000000000000000", "000011110000000", "000000000001111", "000110010100111", "000000000000000", "000000110011111", "000000000000000", "000000010100011", "000000000000000", "100000111010000", "000000000011110", "000100100101100", "000001001111010", "000000000000000", "000010101001001", "000100011100101", "000010010001011", "100000101010000", "000001100111110", "100000100000111", "000010011011011", "001000110010010", "000000000000000", "100101010110101", "000010100100110", "001001001011111", "100000101001111", "100101111111110", "000000110110101", "100011100001010", "000000001011001", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000000000001010", "101001010100100", "000101000100000", "000001110110111", "000000000000000", "000000010111110", "000000000000000", "000000000000000", "000010111110100", "100001001110001", "000000001001000", "000010101110101", "100001000100000", "110011100010011", "000010110011011", "100000110100011", "000000000000000", "101100101001101", "000011010001111", "100011100000010", "000000000101111", "000100001100110", "000000010000001", "000100111100001", "100000101000010", "000000000000000", "000000000000000", "100001000100101", "000010010001111", "000000000000000", "000000100100011", "000010010100110", "000001111000110", "100001001110010", "000000010111111", "000010110101110", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "000010000011100", "000010111100100", "000000000000000", "000000000000000", "000001000110011", "000000010000000", "000000110110110", "001110111111010", "100001001000110", "100101110101100", "000001011010101", "100100010010001", "000000110011101", "000000011110111", "000000000000000", "100010110000101", "000000010101000", "000000010101110", "000001011110010", "000111000101100", "000000000000000", "101000100010011", "000001001010111", "100101010111101", "000000101110010", "000000011010000", "000000000000000", "100101101010100", "000010000001101", "000000000000000", "000001101011011", "000000000000000", "000010001000111", "000000000001011", "000000000000000", "000001001110000", "000000010110010", "001100000110000", "100000111100100", "000101110011100", "000000000000000", "000000000000000", "000010011011010", "000110001101011", "000000000000000", "000001111101110", "000000000000000", "000000101111000", "000000000000000", "000010001111011", "000000000000000", "100000100101110", "000001100011101", "000001101011100", "000000010100101", "000000000000000", "000001100000011", "000000000000000", "000010100110110", "000101011001011", "000000000000000", "100011101110010", "000011110110010", "000101011001100", "000000011100101", "000100100000100", "000000000000000", "000010010001111", "000000000000000", "100010011011000", "000100011001010", "000000001010010", "000000110100111", "101011011001100", "000010000110011", "100111100001001", "000100000111000", "000000000000000", "000000000000000", "000111111100111", "000000000000000", "100100101101110", "000001011011111", "100011011111001", "000000010100100", "100010001100000", "000000101100010", "100010110100111", "000011101101010", "101100001000110", "000010000100001", "100101010101111", "000001101011100", "000000000000000", "000000111111011", "000000000000000", "000000000000000", "100001000011000", "000001000100100", "000000000000000", "000000000101001", "000001001100101", "000010101100001", "000010101010001", "000000011110100", "000000110000100", "000000011001000", "000001011111110", "000011101111001", "000000000000000", "000010000011100", "001001001000011", "000000000000000", "000100001100110", "000000000000000", "000111100010100", "000000000000000", "000001101100000", "000010010110011", "000101101001100", "000000000000000", "000000010001001", "000000100111100", "000010001111010", "000000000000000", "000010010111101", "000001111111000", "000000000000000", "000000000000000", "100100011001001", "000001101111101", "000000000000000", "000000001101011", "000000000000000", "000000000000000", "100110011100110", "000010011000001", "100111100111111", "000001100011111", "000010010001000", "000000000000000", "000000001111100", "000000000011011", "100000111110011", "000001001100101", "100010100001000", "000010101000011", "100011010110110", "000010101101111", "000010111101101", "000000000000000", "000000000000000", "000000100011110", "000000000000000", "000000000000000", "000010111111010", "000000000000000", "000011100011101", "000001101110010", "000011110000110", "000010101100110", "000011110110110", "000010001001100", "000010110000001", "000001001111111", "000101000010100", "000001010000011", "000000000000000", "000010011010111", "000100011100011", "000000000000000", "000000000000000", "000011010111100", "000000000000000", "000010100001110", "100000100000000", "000010101100001", "100100101110111", "000010110010010", "000100010001111", "000000000000000", "000010000111001", "000000000000000", "000111111001011", "000000000000000", "001010000101110", "000000000000000", "000100011110001", "000000111100101", "100001110001000", "000010001001100", "000010001110011", "000000110111110", "000001111111101", "000000000000000", "100000111001110", "000000000000000", "100001100000111", "000000001100011", "100001000100101", "000000000000000", "000000011000000", "000000000000000", "000001100100010", "000000000000000", "000010110000001", "000000011110001", "000000100110011", "000000000000000", "001000110011011", "100001000100000", "000000100111111", "000001110000000", "000011101000110", "000000100011110", "000000101001011", "000001101100000", "000000000110111", "000010101010001", "000011011011100", "000000101010101", "000011111100111", "000001010000000", "000000011010010", "000011000001011", "000010000101001", "000000000000000", "000000000000000", "000000100001110", "000000000000000", "000010101101100", "000000000100001", "000000000000000", "000000100010010", "000000000000000", "100001111010100", "000000100101010", "100010001011000", "000000101001101", "000000000000000", "000010110011000", "100000101010010", "000000111101100", "000000000000000", "000000000000000", "000001000111000", "000010011111000", "000000000000000", "000000000000000", "000000000000000", "000001100001100", "000000000000000", "000001000101111", "000111111011111", "000000000000000", "000000000000000", "000000000000000", "100100010001100", "000001000101101", "000000000000000", "000010011111100", "000000000000000", "000000000000000", "001001100111110", "000000000000000", "000000010111101", "000000000000000", "000010101011110", "000100111110100", "000100011111010", "000100111100010", "000011111000100", "000001011001100", "000001111111000", "000100010001011", "000100101001001", "000010010000010", "000010010111011", "000011100111101", "000001011110111", "000001111100101", "000010101010011", "000000000110110", "000011000001111", "000000101001111", "000000000000000", "000010010000101", "000001101110010", "000100111100011", "000000000000001", "000001101001011", "100000111010011", "000000011111000", "100001000101100", "000011110011001", "000000010011101", "000010010000110", "000000000000000", "000000000000000", "000000000000000", "000000000000000", "100001110100001", "000001010011111", "000000011001100", "000000101100001", "000000000000000", "000001000011111", "000000000000000", "000010001000100", "000101011100110", "000000000111001", "000010010110001", "000000000000000", "000010010001000", "000000000000000", "000001001100000", "000010101011001", "100010000010101", "000001100101111", "000000110100111", "000000000000000", "000000110101101", "000010000011011", "000000110111000", "000010010110101", "000010011010010", "000100100101110", "000001101100100", "000100000010100", "000000010000010", "000001010110101", "000011000000100", "000001000000000", "000010100111110", "000011101011010", "000010111000110", "000011011100101", "000000100101101", "000100010000101", "000011110001001", "000010000101000", "000011011100100", "000000100100100", "000000000000000", "000000000000000", "000000000000000", "000001111100010", "000010111011110", "000000001110000", "000011100111010", "000100010010000", "000100110000110", "000001010100111", "000000000000000", "000000000000000", "100001101000001", "000000011100001", "100000101101110", "000000000110100", "000000001100100", "000001000011000", "000000000000000", "000000000000000", "100001000100011", "000000100010101", "100010000010101", "000001011111001", "100010000010101", "000010010011000", "100010000010101", "000011010001011", "100001011100001", "000000010101100", "000010110100001", "000001100011100", "000010100110100", "000000100100100", "000010110001000", "000000000000000", "000100101010010", "000000000000000", "000010000001110", "000011110011000", "000100110001110", "000010001011011", "100101100011101", "000001110111101"); 

testO<=test;
layerO<=layer;
process(selecttest,test)
begin
	if selecttest="00" then
		test<= ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0');
		--circle
	elsif selecttest="01" then
		test<= ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0');
		--square
	elsif selecttest="10" then 
		test<= ('0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '1', '1', '1', '1', '1', '1', '1', '1', '1', '1', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0', '0');
		--triangle
	end if;
end process;

process(reset,clk)
variable i : integer range 0 to 784:=0;
	begin 
	if(reset = '1') then
		i:=0;
		state<="00";
		layer		<=((others=> (others=>'0')));
		outputSum<=(others=>'0');
		outputSignal<='0';
	elsif(rising_edge(clk)) then
		case state is 
			when "00"=>
				if i<=783 then
					layer(0)<=sum1815(x=>layer(0),y=>mulIw1(I=>test(i),w1=>weight(i*2)));
					layer(1)<=sum1815(x=>layer(1),y=>mulIw1(I=>test(i),w1=>weight(i*2+1)));
					i:=i+1;
				else	
					layer(0)<=sigmoid18(layer(0));
					layer(1)<=sigmoid18(layer(1));
					state <="01";
				end if;
			when "01"=>
				outputSum<=sum1515(x=>mullw2(	l1=>layer(0),w2=>weight(1568)	),y=>mullw2(l1=>layer(1),w2=>weight(1569)));
				state <="10";
			when "10"=>
			outputSum<=sigmoid18(outputSum);
			state<="11";
			when others=>
			outputSignal<=(outputSum(8) or outputSum(7));
		end case;
	end if;
end process;

end rtl;
