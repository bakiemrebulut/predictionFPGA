LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.ALL;


ENTITY hw_image_generator IS
  PORT(
		ready	 :	 IN 	std_logic;
		clk		: in std_logic;
		dataIn	 :	 IN 	std_logic_vector(0 downto 0);
		address	 :	 out	STD_LOGIC_VECTOR(16 DOWNTO 0);

		disp_ena :	IN	STD_LOGIC;
		row      :  IN   INTEGER;    --row pixel coordinate
		column   :  IN   INTEGER;    --column pixel coordinate
		screenEnable: IN std_logic;
		annout	:  IN std_LOGIC;
		red      :  OUT  STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => '0');  --red magnitude output to DAC
		green    :  OUT  STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => '0');  --green magnitude output to DAC
		blue     :  OUT  STD_LOGIC_VECTOR(0 DOWNTO 0) := (OTHERS => '0')); --blue magnitude output to DAC
END hw_image_generator;

ARCHITECTURE behavior OF hw_image_generator IS

signal redS   : std_logic_vector(0 downto 0);
signal greenS : std_logic_vector(0 downto 0);
signal blueS  : std_logic_vector(0 downto 0);
signal addressSignal:std_LOGIC_VECTOR(16 DOWNTO 0);
signal annrate : integer range 0 to 997:=0;
signal scrEnLatch : std_logic;
type rom_type is array (0 to 159 , 0 to 7) of std_logic_vector(0 downto 0);
signal ROM: rom_type := (("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","1","1","1","1","1","0","0"),("1","1","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("1","1","0","0","1","1","1","0"),("1","1","0","1","1","1","1","0"),("1","1","1","1","0","1","1","0"),("1","1","1","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("0","1","1","1","1","1","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","1","1","0","0","0"),("0","0","1","1","1","0","0","0"),("0","1","1","1","1","0","0","0"),("0","0","0","1","1","0","0","0"),("0","0","0","1","1","0","0","0"),("0","0","0","1","1","0","0","0"),("0","0","0","1","1","0","0","0"),("0","0","0","1","1","0","0","0"),("0","0","0","1","1","0","0","0"),("0","1","1","1","1","1","1","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","1","1","1","1","1","0","0"),("1","1","0","0","0","1","1","0"),("0","0","0","0","0","1","1","0"),("0","0","0","0","1","1","0","0"),("0","0","0","1","1","0","0","0"),("0","0","1","1","0","0","0","0"),("0","1","1","0","0","0","0","0"),("1","1","0","0","0","0","0","0"),("1","1","0","0","0","1","1","0"),("1","1","1","1","1","1","1","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","1","1","1","1","1","0","0"),("1","1","0","0","0","1","1","0"),("0","0","0","0","0","1","1","0"),("0","0","0","0","0","1","1","0"),("0","0","1","1","1","1","0","0"),("0","0","0","0","0","1","1","0"),("0","0","0","0","0","1","1","0"),("0","0","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("0","1","1","1","1","1","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","1","1","0","0"),("0","0","0","1","1","1","0","0"),("0","0","1","1","1","1","0","0"),("0","1","1","0","1","1","0","0"),("1","1","0","0","1","1","0","0"),("1","1","1","1","1","1","1","0"),("0","0","0","0","1","1","0","0"),("0","0","0","0","1","1","0","0"),("0","0","0","0","1","1","0","0"),("0","0","0","1","1","1","1","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("1","1","1","1","1","1","1","0"),("1","1","0","0","0","0","0","0"),("1","1","0","0","0","0","0","0"),("1","1","0","0","0","0","0","0"),("1","1","1","1","1","1","0","0"),("0","0","0","0","0","1","1","0"),("0","0","0","0","0","1","1","0"),("0","0","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("0","1","1","1","1","1","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","1","1","1","0","0","0"),("0","1","1","0","0","0","0","0"),("1","1","0","0","0","0","0","0"),("1","1","0","0","0","0","0","0"),("1","1","1","1","1","1","0","0"),("1","1","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("0","1","1","1","1","1","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("1","1","1","1","1","1","1","0"),("1","1","0","0","0","1","1","0"),("0","0","0","0","0","1","1","0"),("0","0","0","0","0","1","1","0"),("0","0","0","0","1","1","0","0"),("0","0","0","1","1","0","0","0"),("0","0","1","1","0","0","0","0"),("0","0","1","1","0","0","0","0"),("0","0","1","1","0","0","0","0"),("0","0","1","1","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","1","1","1","1","1","0","0"),("1","1","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("0","1","1","1","1","1","0","0"),("1","1","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("0","1","1","1","1","1","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","1","1","1","1","1","0","0"),("1","1","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("1","1","0","0","0","1","1","0"),("0","1","1","1","1","1","1","0"),("0","0","0","0","0","1","1","0"),("0","0","0","0","0","1","1","0"),("0","0","0","0","0","1","1","0"),("0","0","0","0","1","1","0","0"),("0","1","1","1","1","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"),("0","0","0","0","0","0","0","0"));
BEGIN
red<=redS;
green<=greenS;
blue<=blueS;
--address<=addressSignal;


PROCESS(clk)
BEGIN
if screenEnable='1' then
	scrEnLatch<=screenEnable;
end if;
address<=std_logic_vector(to_unsigned(row*320+column,addressSignal'length));
if row<=240 and column<=320  then
	if (row=0 or row=240 or column=0 or column=320) then --or((row<232 and row>8 and (column=48 or column=272)) or ((row=8 or row=232) and column>48 and column<272))then
		redS<="1";
		greenS<="1";
		blueS<="1";
		elsif scrEnLatch='1' and screenEnable='1' then
			redS<=dataIn;
			greenS<=dataIn;
			blueS<=dataIn;	
		else 
			redS<="0";
			greenS<="0";
			blueS<="0";
--	else 
--		redS<=dataIn;
--		greenS<=dataIn;
--		blueS<=dataIn;
	end if;
elsif (row>106 and row<135) and (column>320 and column<349) then
	address<=std_logic_vector(to_unsigned(76800+(row-107)*28+(column-321),addressSignal'length));
	redS<=dataIn;
	greenS<=dataIn;
	blueS<=dataIn;
elsif (row>112 and row<112+16*2+1) and (column>350 and column<350+8*2+1) then--d1
	if annout='0' then
		redS<=ROM((row-113)/2,(column-351)/2);
		greenS<="0";
		blueS<="0";
	else
		redS<=ROM((row-113)/2+16,(column-351)/2);
		greenS<="0";
		blueS<="0";
	end if;

else
	redS<="0";
	greenS<="0";
	blueS<="0";
end if;

end process;
END behavior;
